
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/21/2024 10:40:22 AM
// Design Name: 
// Module Name: intmul32_64_top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module intmul(input clk,rst,
              input [254:0] A,
              input [254:0] B,
              output reg [509:0] D);


(* use_dsp = "yes" *) reg [40:0] p0_0,p0_1,p0_2,p0_3,p0_4,p0_5,p0_6,p0_7,p0_8,p0_9,p0_10,p1_0,p1_1,p1_2,p1_3,p1_4,p1_5,p1_6,p1_7,p1_8,p1_9,p1_10,p2_0,p2_1,p2_2,p2_3,p2_4,p2_5,p2_6,p2_7,p2_8,p2_9,p2_10,p3_0,p3_1,p3_2,p3_3,p3_4,p3_5,p3_6,p3_7,p3_8,p3_9,p3_10,p4_0,p4_1,p4_2,p4_3,p4_4,p4_5,p4_6,p4_7,p4_8,p4_9,p4_10,p5_0,p5_1,p5_2,p5_3,p5_4,p5_5,p5_6,p5_7,p5_8,p5_9,p5_10,p6_0,p6_1,p6_2,p6_3,p6_4,p6_5,p6_6,p6_7,p6_8,p6_9,p6_10,p7_0,p7_1,p7_2,p7_3,p7_4,p7_5,p7_6,p7_7,p7_8,p7_9,p7_10,p8_0,p8_1,p8_2,p8_3,p8_4,p8_5,p8_6,p8_7,p8_8,p8_9,p8_10,p9_0,p9_1,p9_2,p9_3,p9_4,p9_5,p9_6,p9_7,p9_8,p9_9,p9_10,p10_0,p10_1,p10_2,p10_3,p10_4,p10_5,p10_6,p10_7,p10_8,p10_9,p10_10,p11_0,p11_1,p11_2,p11_3,p11_4,p11_5,p11_6,p11_7,p11_8,p11_9,p11_10,p12_0,p12_1,p12_2,p12_3,p12_4,p12_5,p12_6,p12_7,p12_8,p12_9,p12_10,p13_0,p13_1,p13_2,p13_3,p13_4,p13_5,p13_6,p13_7,p13_8,p13_9,p13_10,p14_0,p14_1,p14_2,p14_3,p14_4,p14_5,p14_6,p14_7,p14_8,p14_9,p14_10;


always @(posedge clk or posedge rst) begin
    if(rst) begin
        p0_0 <= 0;
        p0_1 <= 0;
        p0_2 <= 0;
        p0_3 <= 0;
        p0_4 <= 0;
        p0_5 <= 0;
        p0_6 <= 0;
        p0_7 <= 0;
        p0_8 <= 0;
        p0_9 <= 0;
        p0_10 <= 0;
        p1_0 <= 0;
        p1_1 <= 0;
        p1_2 <= 0;
        p1_3 <= 0;
        p1_4 <= 0;
        p1_5 <= 0;
        p1_6 <= 0;
        p1_7 <= 0;
        p1_8 <= 0;
        p1_9 <= 0;
        p1_10 <= 0;
        p2_0 <= 0;
        p2_1 <= 0;
        p2_2 <= 0;
        p2_3 <= 0;
        p2_4 <= 0;
        p2_5 <= 0;
        p2_6 <= 0;
        p2_7 <= 0;
        p2_8 <= 0;
        p2_9 <= 0;
        p2_10 <= 0;
        p3_0 <= 0;
        p3_1 <= 0;
        p3_2 <= 0;
        p3_3 <= 0;
        p3_4 <= 0;
        p3_5 <= 0;
        p3_6 <= 0;
        p3_7 <= 0;
        p3_8 <= 0;
        p3_9 <= 0;
        p3_10 <= 0;
        p4_0 <= 0;
        p4_1 <= 0;
        p4_2 <= 0;
        p4_3 <= 0;
        p4_4 <= 0;
        p4_5 <= 0;
        p4_6 <= 0;
        p4_7 <= 0;
        p4_8 <= 0;
        p4_9 <= 0;
        p4_10 <= 0;
        p5_0 <= 0;
        p5_1 <= 0;
        p5_2 <= 0;
        p5_3 <= 0;
        p5_4 <= 0;
        p5_5 <= 0;
        p5_6 <= 0;
        p5_7 <= 0;
        p5_8 <= 0;
        p5_9 <= 0;
        p5_10 <= 0;
        p6_0 <= 0;
        p6_1 <= 0;
        p6_2 <= 0;
        p6_3 <= 0;
        p6_4 <= 0;
        p6_5 <= 0;
        p6_6 <= 0;
        p6_7 <= 0;
        p6_8 <= 0;
        p6_9 <= 0;
        p6_10 <= 0;
        p7_0 <= 0;
        p7_1 <= 0;
        p7_2 <= 0;
        p7_3 <= 0;
        p7_4 <= 0;
        p7_5 <= 0;
        p7_6 <= 0;
        p7_7 <= 0;
        p7_8 <= 0;
        p7_9 <= 0;
        p7_10 <= 0;
        p8_0 <= 0;
        p8_1 <= 0;
        p8_2 <= 0;
        p8_3 <= 0;
        p8_4 <= 0;
        p8_5 <= 0;
        p8_6 <= 0;
        p8_7 <= 0;
        p8_8 <= 0;
        p8_9 <= 0;
        p8_10 <= 0;
        p9_0 <= 0;
        p9_1 <= 0;
        p9_2 <= 0;
        p9_3 <= 0;
        p9_4 <= 0;
        p9_5 <= 0;
        p9_6 <= 0;
        p9_7 <= 0;
        p9_8 <= 0;
        p9_9 <= 0;
        p9_10 <= 0;
        p10_0 <= 0;
        p10_1 <= 0;
        p10_2 <= 0;
        p10_3 <= 0;
        p10_4 <= 0;
        p10_5 <= 0;
        p10_6 <= 0;
        p10_7 <= 0;
        p10_8 <= 0;
        p10_9 <= 0;
        p10_10 <= 0;
        p11_0 <= 0;
        p11_1 <= 0;
        p11_2 <= 0;
        p11_3 <= 0;
        p11_4 <= 0;
        p11_5 <= 0;
        p11_6 <= 0;
        p11_7 <= 0;
        p11_8 <= 0;
        p11_9 <= 0;
        p11_10 <= 0;
        p12_0 <= 0;
        p12_1 <= 0;
        p12_2 <= 0;
        p12_3 <= 0;
        p12_4 <= 0;
        p12_5 <= 0;
        p12_6 <= 0;
        p12_7 <= 0;
        p12_8 <= 0;
        p12_9 <= 0;
        p12_10 <= 0;
        p13_0 <= 0;
        p13_1 <= 0;
        p13_2 <= 0;
        p13_3 <= 0;
        p13_4 <= 0;
        p13_5 <= 0;
        p13_6 <= 0;
        p13_7 <= 0;
        p13_8 <= 0;
        p13_9 <= 0;
        p13_10 <= 0;
        p14_0 <= 0;
        p14_1 <= 0;
        p14_2 <= 0;
        p14_3 <= 0;
        p14_4 <= 0;
        p14_5 <= 0;
        p14_6 <= 0;
        p14_7 <= 0;
        p14_8 <= 0;
        p14_9 <= 0;
        p14_10 <= 0;


    end
    else begin
        p0_0 <= A[16:0] * B[23:0];
        p0_1 <= A[16:0] * B[47:24];
        p0_2 <= A[16:0] * B[71:48];
        p0_3 <= A[16:0] * B[95:72];
        p0_4 <= A[16:0] * B[119:96];
        p0_5 <= A[16:0] * B[143:120];
        p0_6 <= A[16:0] * B[167:144];
        p0_7 <= A[16:0] * B[191:168];
        p0_8 <= A[16:0] * B[215:192];
        p0_9 <= A[16:0] * B[239:216];
        p0_10 <= A[16:0] * B[254:240];
        p1_0 <= A[33:17] * B[23:0];
        p1_1 <= A[33:17] * B[47:24];
        p1_2 <= A[33:17] * B[71:48];
        p1_3 <= A[33:17] * B[95:72];
        p1_4 <= A[33:17] * B[119:96];
        p1_5 <= A[33:17] * B[143:120];
        p1_6 <= A[33:17] * B[167:144];
        p1_7 <= A[33:17] * B[191:168];
        p1_8 <= A[33:17] * B[215:192];
        p1_9 <= A[33:17] * B[239:216];
        p1_10 <= A[33:17] * B[254:240];
        p2_0 <= A[50:34] * B[23:0];
        p2_1 <= A[50:34] * B[47:24];
        p2_2 <= A[50:34] * B[71:48];
        p2_3 <= A[50:34] * B[95:72];
        p2_4 <= A[50:34] * B[119:96];
        p2_5 <= A[50:34] * B[143:120];
        p2_6 <= A[50:34] * B[167:144];
        p2_7 <= A[50:34] * B[191:168];
        p2_8 <= A[50:34] * B[215:192];
        p2_9 <= A[50:34] * B[239:216];
        p2_10 <= A[50:34] * B[254:240];
        p3_0 <= A[67:51] * B[23:0];
        p3_1 <= A[67:51] * B[47:24];
        p3_2 <= A[67:51] * B[71:48];
        p3_3 <= A[67:51] * B[95:72];
        p3_4 <= A[67:51] * B[119:96];
        p3_5 <= A[67:51] * B[143:120];
        p3_6 <= A[67:51] * B[167:144];
        p3_7 <= A[67:51] * B[191:168];
        p3_8 <= A[67:51] * B[215:192];
        p3_9 <= A[67:51] * B[239:216];
        p3_10 <= A[67:51] * B[254:240];
        p4_0 <= A[84:68] * B[23:0];
        p4_1 <= A[84:68] * B[47:24];
        p4_2 <= A[84:68] * B[71:48];
        p4_3 <= A[84:68] * B[95:72];
        p4_4 <= A[84:68] * B[119:96];
        p4_5 <= A[84:68] * B[143:120];
        p4_6 <= A[84:68] * B[167:144];
        p4_7 <= A[84:68] * B[191:168];
        p4_8 <= A[84:68] * B[215:192];
        p4_9 <= A[84:68] * B[239:216];
        p4_10 <= A[84:68] * B[254:240];
        p5_0 <= A[101:85] * B[23:0];
        p5_1 <= A[101:85] * B[47:24];
        p5_2 <= A[101:85] * B[71:48];
        p5_3 <= A[101:85] * B[95:72];
        p5_4 <= A[101:85] * B[119:96];
        p5_5 <= A[101:85] * B[143:120];
        p5_6 <= A[101:85] * B[167:144];
        p5_7 <= A[101:85] * B[191:168];
        p5_8 <= A[101:85] * B[215:192];
        p5_9 <= A[101:85] * B[239:216];
        p5_10 <= A[101:85] * B[254:240];
        p6_0 <= A[118:102] * B[23:0];
        p6_1 <= A[118:102] * B[47:24];
        p6_2 <= A[118:102] * B[71:48];
        p6_3 <= A[118:102] * B[95:72];
        p6_4 <= A[118:102] * B[119:96];
        p6_5 <= A[118:102] * B[143:120];
        p6_6 <= A[118:102] * B[167:144];
        p6_7 <= A[118:102] * B[191:168];
        p6_8 <= A[118:102] * B[215:192];
        p6_9 <= A[118:102] * B[239:216];
        p6_10 <= A[118:102] * B[254:240];
        p7_0 <= A[135:119] * B[23:0];
        p7_1 <= A[135:119] * B[47:24];
        p7_2 <= A[135:119] * B[71:48];
        p7_3 <= A[135:119] * B[95:72];
        p7_4 <= A[135:119] * B[119:96];
        p7_5 <= A[135:119] * B[143:120];
        p7_6 <= A[135:119] * B[167:144];
        p7_7 <= A[135:119] * B[191:168];
        p7_8 <= A[135:119] * B[215:192];
        p7_9 <= A[135:119] * B[239:216];
        p7_10 <= A[135:119] * B[254:240];
        p8_0 <= A[152:136] * B[23:0];
        p8_1 <= A[152:136] * B[47:24];
        p8_2 <= A[152:136] * B[71:48];
        p8_3 <= A[152:136] * B[95:72];
        p8_4 <= A[152:136] * B[119:96];
        p8_5 <= A[152:136] * B[143:120];
        p8_6 <= A[152:136] * B[167:144];
        p8_7 <= A[152:136] * B[191:168];
        p8_8 <= A[152:136] * B[215:192];
        p8_9 <= A[152:136] * B[239:216];
        p8_10 <= A[152:136] * B[254:240];
        p9_0 <= A[169:153] * B[23:0];
        p9_1 <= A[169:153] * B[47:24];
        p9_2 <= A[169:153] * B[71:48];
        p9_3 <= A[169:153] * B[95:72];
        p9_4 <= A[169:153] * B[119:96];
        p9_5 <= A[169:153] * B[143:120];
        p9_6 <= A[169:153] * B[167:144];
        p9_7 <= A[169:153] * B[191:168];
        p9_8 <= A[169:153] * B[215:192];
        p9_9 <= A[169:153] * B[239:216];
        p9_10 <= A[169:153] * B[254:240];
        p10_0 <= A[186:170] * B[23:0];
        p10_1 <= A[186:170] * B[47:24];
        p10_2 <= A[186:170] * B[71:48];
        p10_3 <= A[186:170] * B[95:72];
        p10_4 <= A[186:170] * B[119:96];
        p10_5 <= A[186:170] * B[143:120];
        p10_6 <= A[186:170] * B[167:144];
        p10_7 <= A[186:170] * B[191:168];
        p10_8 <= A[186:170] * B[215:192];
        p10_9 <= A[186:170] * B[239:216];
        p10_10 <= A[186:170] * B[254:240];
        p11_0 <= A[203:187] * B[23:0];
        p11_1 <= A[203:187] * B[47:24];
        p11_2 <= A[203:187] * B[71:48];
        p11_3 <= A[203:187] * B[95:72];
        p11_4 <= A[203:187] * B[119:96];
        p11_5 <= A[203:187] * B[143:120];
        p11_6 <= A[203:187] * B[167:144];
        p11_7 <= A[203:187] * B[191:168];
        p11_8 <= A[203:187] * B[215:192];
        p11_9 <= A[203:187] * B[239:216];
        p11_10 <= A[203:187] * B[254:240];
        p12_0 <= A[220:204] * B[23:0];
        p12_1 <= A[220:204] * B[47:24];
        p12_2 <= A[220:204] * B[71:48];
        p12_3 <= A[220:204] * B[95:72];
        p12_4 <= A[220:204] * B[119:96];
        p12_5 <= A[220:204] * B[143:120];
        p12_6 <= A[220:204] * B[167:144];
        p12_7 <= A[220:204] * B[191:168];
        p12_8 <= A[220:204] * B[215:192];
        p12_9 <= A[220:204] * B[239:216];
        p12_10 <= A[220:204] * B[254:240];
        p13_0 <= A[237:221] * B[23:0];
        p13_1 <= A[237:221] * B[47:24];
        p13_2 <= A[237:221] * B[71:48];
        p13_3 <= A[237:221] * B[95:72];
        p13_4 <= A[237:221] * B[119:96];
        p13_5 <= A[237:221] * B[143:120];
        p13_6 <= A[237:221] * B[167:144];
        p13_7 <= A[237:221] * B[191:168];
        p13_8 <= A[237:221] * B[215:192];
        p13_9 <= A[237:221] * B[239:216];
        p13_10 <= A[237:221] * B[254:240];
        p14_0 <= A[254:238] * B[23:0];
        p14_1 <= A[254:238] * B[47:24];
        p14_2 <= A[254:238] * B[71:48];
        p14_3 <= A[254:238] * B[95:72];
        p14_4 <= A[254:238] * B[119:96];
        p14_5 <= A[254:238] * B[143:120];
        p14_6 <= A[254:238] * B[167:144];
        p14_7 <= A[254:238] * B[191:168];
        p14_8 <= A[254:238] * B[215:192];
        p14_9 <= A[254:238] * B[239:216];
        p14_10 <= A[254:238] * B[254:240];

    end
end

wire [509:0] p;



assign p = {{68'b0,p10_10,p9_9,p8_8,p7_7,p6_6,p5_5,p4_4,p3_3,p2_2,p1_1,p0_0}} + {{85'b0,p9_10,p8_9,p7_8,p6_7,p5_6,p4_5,p3_4,p2_3,p1_2,p0_1,24'b0}} + {{102'b0,p8_10,p7_9,p6_8,p5_7,p4_6,p3_5,p2_4,p1_3,p0_2,48'b0}} + {{119'b0,p7_10,p6_9,p5_8,p4_7,p3_6,p2_5,p1_4,p0_3,72'b0}} + {{136'b0,p6_10,p5_9,p4_8,p3_7,p2_6,p1_5,p0_4,96'b0}} + {{153'b0,p5_10,p4_9,p3_8,p2_7,p1_6,p0_5,120'b0}} + {{170'b0,p4_10,p3_9,p2_8,p1_7,p0_6,144'b0}} + {{187'b0,p3_10,p2_9,p1_8,p0_7,168'b0}} + {{204'b0,p2_10,p1_9,p0_8,192'b0}} + {{221'b0,p1_10,p0_9,216'b0}} + {{238'b0,p0_10,240'b0}} + {{51'b0,p11_10,p10_9,p9_8,p8_7,p7_6,p6_5,p5_4,p4_3,p3_2,p2_1,p1_0,17'b0}} + {{34'b0,p12_10,p11_9,p10_8,p9_7,p8_6,p7_5,p6_4,p5_3,p4_2,p3_1,p2_0,34'b0}} + {{17'b0,p13_10,p12_9,p11_8,p10_7,p9_6,p8_5,p7_4,p6_3,p5_2,p4_1,p3_0,51'b0}} + {{p14_10,p13_9,p12_8,p11_7,p10_6,p9_5,p8_4,p7_3,p6_2,p5_1,p4_0,68'b0}} + {{15'b0,p14_9,p13_8,p12_7,p11_6,p10_5,p9_4,p8_3,p7_2,p6_1,p5_0,85'b0}} + {{39'b0,p14_8,p13_7,p12_6,p11_5,p10_4,p9_3,p8_2,p7_1,p6_0,102'b0}} + {{63'b0,p14_7,p13_6,p12_5,p11_4,p10_3,p9_2,p8_1,p7_0,119'b0}} + {{87'b0,p14_6,p13_5,p12_4,p11_3,p10_2,p9_1,p8_0,136'b0}} + {{111'b0,p14_5,p13_4,p12_3,p11_2,p10_1,p9_0,153'b0}} + {{135'b0,p14_4,p13_3,p12_2,p11_1,p10_0,170'b0}} + {{159'b0,p14_3,p13_2,p12_1,p11_0,187'b0}} + {{183'b0,p14_2,p13_1,p12_0,204'b0}} + {{207'b0,p14_1,p13_0,221'b0}} + {{231'b0,p14_0,238'b0}}; 


always @(posedge clk) begin
    D <= p;
end
          
endmodule


